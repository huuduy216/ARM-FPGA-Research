module notGate(in,out);
	input wire in;
	output wire out;
	assign out = !in;
endmodule 