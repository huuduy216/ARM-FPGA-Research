module top();

cpu cpu1();

endmodule