module instMem(input [31:0]progCount, output reg [31:0]inst);
	reg [31:0]instructions[15:0];

	initial begin
	instructions[0] = 32'b10010001000000011011111111100001; //addi X1, X31, 111
	instructions[1] = 32'b10010001000000000101101111100010; //addi X2, X31, 22
	instructions[2] = 32'b10010001000000001000011111100011; //addi X3, X31, 33
	instructions[3] = 32'b10010001000000010011001111100100; //addi X4, X31, 76
	instructions[4] = 32'b10001011000000110000000001000101; //add X5, X5, X3
	instructions[5] = 32'b11010001000000001101110000100110; //subi X6, X1, 55
	instructions[6] = 32'b11001011000000100000000010000111; //sub X7, X4, X2
	instructions[7] = 32'b11111000010000000000000011101000; //ldur X8, [X7, 0];
	instructions[8] = 32'b10001010000001110000000100001001; //and X9, X8, X7
	instructions[9] = 32'b10101010000111110000001111101010; //orr X10, X31, X31
	instructions[10] = 32'b11111000000000000000000000101011; //stur X11, [X1, 0]
	instructions[11] = 32'b10010001000000000001001111101100; //addi X12, X31, 4
	instructions[12] = 32'b11010001000000000000010110001100; //subi X12, X12, 1
	instructions[13] = 32'b10110101000000000000000110001100; //cbnz X12, 12
	instructions[14] = 32'b11111000000001100100001111100111; //stur X7, [X31, 100]
	instructions[15] = 32'b10010001000000010001011111111011; //addi X27, X31, 69
	end
	always @ * begin
	#1 inst = instructions[progCount + 1];
	
	end
endmodule